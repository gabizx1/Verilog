module driver7seg (
   input [3:0] b, 
	output [6:0] d;
);
	
always @ 
begin 
	case (b)
			//numeros
			4'b0000: d = 7'b0111111; 
			4'b0001: d = 7'b0000110; 
			4'b0010: d = 7'b1011011; 
			4'b0011: d = 7'b1001111; 
			4'b0100: d = 7'b1100110; 
			4'b0101: d = 7'b1101101; 
			4'b0110: d = 7'b1111101; 
			4'b0111: d = 7'b0000111; 
			4'b1000: d = 7'b1111111; 
			4'b1001: d = 7'b1101111;
			//letras
			4'b1010: d = 7'b1110111;
			4'b1011: d = 7'b1111100;
			4'b1100: d = 7'b0111001;
			4'b1101: d = 7'b1011110;
			4'b1110: d = 7'b1111001;
			4'b1111: d = 7'b1110001;
			//default: d= 7'b1111111;
	endcase
end

endmodule